Primer disseny Custom (cada transistor és dissenyat)
.include mosfet.model

*Capacitat residual dels transistors
*CL vo GND 1p
*INPUTS
VCfont Vc GND pulse(0 5V 0s 1ps 1ps 10ns 20ns)
VBfont Vb GND pulse(0 5V 0s 1ps 1ps 20ns 40ns)
VAfont Va GND pulse(0 5v 0s 1ps 1ps 40ns 80ns)

*VDD Supply voltage
vddfont Vdd GND dc 5V

*Circuit TRANSISTORS
*VA Inverter
MPA 1 Va Vdd Vdd pfet W=3u L=2u
MNA 1 Va GND GND nfet W=3u L=2u

*PMOS of F = A' + B' * C'

MPNA Vf 1 Vdd Vdd pfet W=3u L=2u
MPB 2 Vb Vdd Vdd pfet W=3u L=2u
MPC Vf Vc 2 Vdd pfet W=3u L=2u

*NMOS of F = (A*(B + C))'

MNNA Vf 1 4 GND nfet W=3u L=2u
MNB 4 Vb GND GND nfet W=3u L=2u
MPC 4 Vc GND GND nfet W=3u L=2u


.tran 20p 80ns 0 40p
*.tran printMostresAlTerminal tempsFinal tempsInical SeparacioEntreMostres

.control
run
plot v(Va)+30 v(Vb)+20 v(Vc)+10 v(2)
plot v(4)

.endc
.end