magic
tech scmos
timestamp 1609148708
<< nwell >>
rect -4 -4 8 6
<< polysilicon >>
rect 1 -1 3 1
rect 1 -8 3 -4
rect -4 -10 3 -8
rect 1 -14 3 -10
rect 1 -19 3 -17
<< ndiffusion >>
rect 0 -17 1 -14
rect 3 -17 4 -14
<< pdiffusion >>
rect 0 -4 1 -1
rect 3 -4 4 -1
<< metal1 >>
rect -4 3 8 6
rect -4 0 0 3
rect 4 -14 8 -4
rect -4 -19 0 -18
<< ntransistor >>
rect 1 -17 3 -14
<< ptransistor >>
rect 1 -4 3 -1
<< ndcontact >>
rect -4 -18 0 -14
rect 4 -18 8 -14
<< pdcontact >>
rect -4 -4 0 0
rect 4 -4 8 0
<< labels >>
rlabel polysilicon -3 -9 -3 -9 3 vA!
rlabel metal1 7 -9 7 -9 7 vnA!
rlabel ndcontact -3 -16 -3 -16 1 GND!
rlabel pdcontact -3 -2 -3 -2 3 Vdd!
<< end >>
