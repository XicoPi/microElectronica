magic
tech scmos
timestamp 1608544210
<< nwell >>
rect -12 -15 13 9
<< polysilicon >>
rect -5 7 -3 9
rect 1 7 3 9
rect 6 7 8 9
rect -5 -5 -3 -4
rect -7 -7 -3 -5
rect -7 -25 -5 -7
rect 1 -25 3 -15
rect 6 -21 8 -15
rect 6 -23 11 -21
rect 9 -25 11 -23
rect -7 -34 -5 -32
rect 1 -34 3 -32
rect 9 -34 11 -32
<< ndiffusion >>
rect -8 -32 -7 -25
rect -5 -32 -4 -25
rect 0 -32 1 -25
rect 3 -28 9 -25
rect 3 -32 4 -28
rect 8 -32 9 -28
rect 11 -32 12 -25
<< pdiffusion >>
rect -8 6 -5 7
rect -6 -4 -5 6
rect -3 -4 1 7
rect -2 -8 1 -4
rect 0 -15 1 -8
rect 3 -15 6 7
rect 8 -15 9 7
<< metal1 >>
rect -12 7 13 9
rect -12 6 9 7
rect -12 -4 -10 6
rect -12 -8 -8 -4
rect -12 -18 0 -15
rect -12 -25 -8 -18
rect -4 -25 16 -22
rect 4 -35 8 -32
rect -12 -36 15 -35
rect -12 -38 4 -36
rect 8 -38 15 -36
<< ntransistor >>
rect -7 -32 -5 -25
rect 1 -32 3 -25
rect 9 -32 11 -25
<< ptransistor >>
rect -5 -4 -3 7
rect 1 -15 3 7
rect 6 -15 8 7
<< ndcontact >>
rect -12 -32 -8 -25
rect -4 -32 0 -25
rect 4 -32 8 -28
rect 12 -32 16 -25
<< pdcontact >>
rect -10 -4 -6 6
rect -4 -15 0 -8
rect 9 -15 13 7
<< psubstratepcontact >>
rect 4 -40 8 -36
<< nsubstratencontact >>
rect -12 -12 -8 -8
<< end >>
