Primer disseny Custom (cada transistor és dissenyat)

*Capacitat residual dels transistors
*CL vo GND 1p
*INPUTS
VCfont Vc GND pulse(0 5V 0s 1ps 1ps 10ns 20ns)
VBfont Vb GND pulse(0 5V 0s 1ps 1ps 20ns 40ns)
VAfont Va GND pulse(0 5v 0s 1ps 1ps 40ns 80ns)

*VDD Supply voltage
vddfont Vdd GND dc 5V

*Circuit TRANSISTORS
*VA Inverter
MNA Vna Va GND GND nfet W=3u L=2u
MPA Vna Va Vdd Vdd pfet W=3u L=2u

*PMOS of F = A' + B' * C'

MPNA Vf Vna Vdd Vdd pfet W=3u L=2u
MPB VcD Vb Vdd Vdd pfet W=3u L=2u
MPC Vf Vc VcD Vdd pfet W=3u L=2u

*NMOS of F = (A*(B + C))'

MNNA Vf Vna Vcbn GND nfet W=3u L=2u
MNB Vnas Vb GND GND nfet W=3u L=2u
MPC Vnas Vc GND GND nfet W=3u L=2u


.tran 20p 80ns 0 40p
*.tran printMostresAlTerminal tempsFinal tempsInical SeparacioEntreMostres

.control
run
plot v(Va)+30 v(Vb)+20 v(Vc)+10 v(Vf)

.endc
.end