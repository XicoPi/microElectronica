* SPICE3 file created from Porta_CMOS.ext - technology: scmos

M1000 vF vnA Vdd Vdd pfet w=13u l=2u
+  ad=99p pd=60u as=201p ps=112u
M1001 Porta_CMOS_part2_0/a_3_n15# vB vF Vdd pfet w=24u l=2u
+  ad=72p pd=54u as=0p ps=0u
M1002 Vdd vC Porta_CMOS_part2_0/a_3_n15# Vdd pfet w=24u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 Porta_CMOS_part2_0/a_n5_n33# vnA GND Gnd nfet w=8u l=2u
+  ad=88p pd=54u as=59p ps=44u
M1004 vF vB Porta_CMOS_part2_0/a_n5_n33# Gnd nfet w=8u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1005 Porta_CMOS_part2_0/a_n5_n33# vC vF Gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1006 vnA vA Vdd Vdd pfet w=3u l=2u
+  ad=19p pd=18u as=0p ps=0u
M1007 vnA vA GND Gnd nfet w=3u l=2u
+  ad=19p pd=18u as=0p ps=0u
C0 Vdd vC 14.58fF
C1 vA GND 14.58fF
C2 Vdd GND 702.14fF
C3 vA Vdd 14.46fF
C4 GND vF 13.50fF
C5 Vdd vF 15.87fF
C6 GND vB 13.50fF
C7 GND vC 13.50fF
C8 Vdd vnA 4.72fF
C9 Vdd vB 14.58fF
C10 vA Gnd 138.14fF
C11 Vdd Gnd 54.98fF
C12 GND Gnd 11.70fF
C13 vF Gnd 6.63fF
C14 vC Gnd 173.46fF
C15 vB Gnd 149.92fF
C16 vnA Gnd 12.62fF
