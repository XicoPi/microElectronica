magic
tech scmos
timestamp 1609168350
<< nwell >>
rect 122 1411 192 1420
rect 122 1408 142 1411
rect 134 1398 142 1408
rect 170 1386 192 1411
<< polysilicon >>
rect 116 1392 122 1394
rect 116 1359 120 1392
rect 136 1385 139 1391
rect 136 1382 142 1385
rect 155 1357 157 1366
rect 163 1357 165 1366
<< metal1 >>
rect 119 1447 163 1448
rect 118 1446 163 1447
rect 117 1445 163 1446
rect 116 1444 163 1445
rect 167 1444 169 1448
rect 173 1444 175 1448
rect 179 1444 181 1448
rect 185 1444 187 1448
rect 191 1447 1405 1448
rect 191 1446 1406 1447
rect 191 1445 1407 1446
rect 191 1444 1408 1445
rect 115 1443 1409 1444
rect 114 1442 1410 1443
rect 113 1441 163 1442
rect 112 1440 163 1441
rect 111 1439 163 1440
rect 110 1438 163 1439
rect 167 1438 169 1442
rect 173 1438 175 1442
rect 179 1438 181 1442
rect 185 1438 187 1442
rect 191 1441 1411 1442
rect 191 1440 1412 1441
rect 191 1439 1413 1440
rect 191 1438 1414 1439
rect 109 1437 121 1438
rect 1403 1437 1415 1438
rect 108 1436 120 1437
rect 1404 1436 1416 1437
rect 107 1435 119 1436
rect 1405 1435 1417 1436
rect 106 1434 118 1435
rect 1406 1434 1418 1435
rect 105 1433 117 1434
rect 1407 1433 1419 1434
rect 104 1432 116 1433
rect 1408 1432 1420 1433
rect 103 1431 115 1432
rect 124 1431 343 1432
rect 102 1430 114 1431
rect 123 1430 343 1431
rect 101 1429 113 1430
rect 122 1429 343 1430
rect 100 1428 112 1429
rect 121 1428 343 1429
rect 347 1428 349 1432
rect 353 1428 355 1432
rect 359 1428 361 1432
rect 365 1428 367 1432
rect 371 1428 433 1432
rect 437 1428 439 1432
rect 443 1428 445 1432
rect 449 1428 451 1432
rect 455 1428 457 1432
rect 461 1428 523 1432
rect 527 1428 529 1432
rect 533 1428 535 1432
rect 539 1428 541 1432
rect 545 1428 547 1432
rect 551 1428 613 1432
rect 617 1428 619 1432
rect 623 1428 625 1432
rect 629 1428 631 1432
rect 635 1428 637 1432
rect 641 1428 703 1432
rect 707 1428 709 1432
rect 713 1428 715 1432
rect 719 1428 721 1432
rect 725 1428 727 1432
rect 731 1428 793 1432
rect 797 1428 799 1432
rect 803 1428 805 1432
rect 809 1428 811 1432
rect 815 1428 817 1432
rect 821 1428 883 1432
rect 887 1428 889 1432
rect 893 1428 895 1432
rect 899 1428 901 1432
rect 905 1428 907 1432
rect 911 1428 973 1432
rect 977 1428 979 1432
rect 983 1428 985 1432
rect 989 1428 991 1432
rect 995 1428 997 1432
rect 1001 1428 1063 1432
rect 1067 1428 1069 1432
rect 1073 1428 1075 1432
rect 1079 1428 1081 1432
rect 1085 1428 1087 1432
rect 1091 1428 1153 1432
rect 1157 1428 1159 1432
rect 1163 1428 1165 1432
rect 1169 1428 1171 1432
rect 1175 1428 1177 1432
rect 1181 1428 1243 1432
rect 1247 1428 1249 1432
rect 1253 1428 1255 1432
rect 1259 1428 1261 1432
rect 1265 1428 1267 1432
rect 1271 1428 1333 1432
rect 1337 1428 1339 1432
rect 1343 1428 1345 1432
rect 1349 1428 1351 1432
rect 1355 1428 1357 1432
rect 1361 1431 1400 1432
rect 1409 1431 1421 1432
rect 1361 1430 1401 1431
rect 1410 1430 1422 1431
rect 1361 1429 1402 1430
rect 1411 1429 1423 1430
rect 1361 1428 1403 1429
rect 1412 1428 1424 1429
rect 99 1427 111 1428
rect 120 1427 1404 1428
rect 1413 1427 1425 1428
rect 98 1426 110 1427
rect 119 1426 1405 1427
rect 1414 1426 1426 1427
rect 97 1425 109 1426
rect 118 1425 343 1426
rect 96 1424 108 1425
rect 117 1424 343 1425
rect 95 1423 107 1424
rect 116 1423 343 1424
rect 94 1422 106 1423
rect 115 1422 343 1423
rect 347 1422 349 1426
rect 353 1422 355 1426
rect 359 1422 361 1426
rect 365 1422 367 1426
rect 371 1422 433 1426
rect 437 1422 439 1426
rect 443 1422 445 1426
rect 449 1422 451 1426
rect 455 1422 457 1426
rect 461 1422 523 1426
rect 527 1422 529 1426
rect 533 1422 535 1426
rect 539 1422 541 1426
rect 545 1422 547 1426
rect 551 1422 613 1426
rect 617 1422 619 1426
rect 623 1422 625 1426
rect 629 1422 631 1426
rect 635 1422 637 1426
rect 641 1422 703 1426
rect 707 1422 709 1426
rect 713 1422 715 1426
rect 719 1422 721 1426
rect 725 1422 727 1426
rect 731 1422 793 1426
rect 797 1422 799 1426
rect 803 1422 805 1426
rect 809 1422 811 1426
rect 815 1422 817 1426
rect 821 1422 883 1426
rect 887 1422 889 1426
rect 893 1422 895 1426
rect 899 1422 901 1426
rect 905 1422 907 1426
rect 911 1422 973 1426
rect 977 1422 979 1426
rect 983 1422 985 1426
rect 989 1422 991 1426
rect 995 1422 997 1426
rect 1001 1422 1063 1426
rect 1067 1422 1069 1426
rect 1073 1422 1075 1426
rect 1079 1422 1081 1426
rect 1085 1422 1087 1426
rect 1091 1422 1153 1426
rect 1157 1422 1159 1426
rect 1163 1422 1165 1426
rect 1169 1422 1171 1426
rect 1175 1422 1177 1426
rect 1181 1422 1243 1426
rect 1247 1422 1249 1426
rect 1253 1422 1255 1426
rect 1259 1422 1261 1426
rect 1265 1422 1267 1426
rect 1271 1422 1333 1426
rect 1337 1422 1339 1426
rect 1343 1422 1345 1426
rect 1349 1422 1351 1426
rect 1355 1422 1357 1426
rect 1361 1425 1406 1426
rect 1415 1425 1427 1426
rect 1361 1424 1407 1425
rect 1416 1424 1428 1425
rect 1361 1423 1408 1424
rect 1417 1423 1429 1424
rect 1361 1422 1409 1423
rect 1418 1422 1430 1423
rect 93 1421 105 1422
rect 114 1421 126 1422
rect 1398 1421 1410 1422
rect 1419 1421 1431 1422
rect 92 1420 104 1421
rect 113 1420 125 1421
rect 1399 1420 1411 1421
rect 1420 1420 1432 1421
rect 91 1419 103 1420
rect 112 1419 124 1420
rect 1400 1419 1412 1420
rect 1421 1419 1433 1420
rect 90 1418 102 1419
rect 111 1418 123 1419
rect 89 1417 101 1418
rect 110 1417 122 1418
rect 88 1416 100 1417
rect 109 1416 121 1417
rect 130 1416 136 1418
rect 87 1415 99 1416
rect 108 1415 120 1416
rect 86 1414 98 1415
rect 107 1414 119 1415
rect 126 1414 136 1416
rect 140 1415 153 1418
rect 1401 1418 1413 1419
rect 1422 1418 1434 1419
rect 157 1415 163 1418
rect 140 1414 163 1415
rect 167 1414 169 1418
rect 173 1414 175 1418
rect 179 1414 181 1418
rect 185 1414 187 1418
rect 191 1414 192 1418
rect 1402 1417 1414 1418
rect 1423 1417 1435 1418
rect 1403 1416 1415 1417
rect 1424 1416 1436 1417
rect 1404 1415 1416 1416
rect 1425 1415 1437 1416
rect 1405 1414 1417 1415
rect 1426 1414 1438 1415
rect 85 1413 97 1414
rect 106 1413 118 1414
rect 124 1413 128 1414
rect 84 1412 96 1413
rect 105 1412 117 1413
rect 123 1412 128 1413
rect 83 1411 95 1412
rect 104 1411 116 1412
rect 82 1410 94 1411
rect 103 1410 115 1411
rect 122 1410 128 1412
rect 132 1411 192 1414
rect 1406 1413 1418 1414
rect 1427 1413 1439 1414
rect 1407 1412 1419 1413
rect 1428 1412 1440 1413
rect 1408 1411 1420 1412
rect 1429 1411 1441 1412
rect 132 1410 142 1411
rect 81 1409 93 1410
rect 102 1409 114 1410
rect 80 1408 92 1409
rect 101 1408 113 1409
rect 122 1408 142 1410
rect 79 1407 91 1408
rect 100 1407 112 1408
rect 78 1406 90 1407
rect 99 1406 111 1407
rect 77 1405 89 1406
rect 98 1405 110 1406
rect 134 1405 142 1408
rect 170 1410 192 1411
rect 1409 1410 1421 1411
rect 1430 1410 1442 1411
rect 76 1404 88 1405
rect 97 1404 109 1405
rect 76 1403 87 1404
rect 96 1403 108 1404
rect 76 121 86 1403
rect 95 1402 107 1403
rect 94 1401 106 1402
rect 93 1400 105 1401
rect 92 1399 104 1400
rect 92 1398 103 1399
rect 92 1379 102 1398
rect 134 1391 135 1395
rect 170 1389 177 1410
rect 1410 1409 1422 1410
rect 1431 1409 1443 1410
rect 1411 1408 1423 1409
rect 1432 1408 1444 1409
rect 1412 1407 1424 1408
rect 1433 1407 1445 1408
rect 1413 1406 1425 1407
rect 1434 1406 1446 1407
rect 1414 1405 1426 1406
rect 1435 1405 1447 1406
rect 1415 1404 1427 1405
rect 1436 1404 1448 1405
rect 1416 1403 1428 1404
rect 1437 1403 1448 1404
rect 1417 1402 1429 1403
rect 1418 1401 1430 1402
rect 1419 1400 1431 1401
rect 1420 1399 1432 1400
rect 1421 1398 1432 1399
rect 122 1379 126 1383
rect 92 1377 129 1379
rect 92 1373 122 1377
rect 126 1376 129 1377
rect 126 1373 142 1376
rect 92 1370 142 1373
rect 92 1091 102 1370
rect 123 1368 142 1370
rect 127 1364 131 1368
rect 135 1366 142 1368
rect 135 1364 146 1366
rect 123 1362 146 1364
rect 109 1360 120 1362
rect 114 1359 120 1360
rect 114 1355 116 1359
rect 109 1352 116 1355
rect 114 1347 116 1352
rect 109 1344 116 1347
rect 114 1339 116 1344
rect 1422 1361 1432 1398
rect 1426 1357 1428 1361
rect 154 1349 158 1353
rect 109 1332 120 1339
rect 123 1345 158 1349
rect 123 1324 128 1345
rect 162 1342 166 1353
rect 109 1319 128 1324
rect 136 1338 166 1342
rect 1422 1355 1432 1357
rect 1426 1351 1428 1355
rect 1422 1349 1432 1351
rect 1426 1345 1428 1349
rect 1422 1343 1432 1345
rect 1426 1339 1428 1343
rect 109 1271 115 1319
rect 136 1314 141 1338
rect 114 1267 115 1271
rect 109 1264 115 1267
rect 114 1260 115 1264
rect 109 1257 115 1260
rect 114 1253 115 1257
rect 109 1250 115 1253
rect 114 1246 115 1250
rect 109 1242 115 1246
rect 120 1310 141 1314
rect 1422 1337 1432 1339
rect 1426 1333 1428 1337
rect 120 1182 124 1310
rect 110 1178 124 1182
rect 110 1174 112 1178
rect 116 1174 119 1178
rect 123 1174 124 1178
rect 110 1171 124 1174
rect 110 1167 112 1171
rect 116 1167 119 1171
rect 123 1167 124 1171
rect 110 1165 124 1167
rect 110 1161 112 1165
rect 116 1161 119 1165
rect 123 1161 124 1165
rect 110 1159 124 1161
rect 110 1155 112 1159
rect 116 1155 119 1159
rect 123 1155 124 1159
rect 110 1152 124 1155
rect 1422 1271 1432 1333
rect 1426 1267 1428 1271
rect 1422 1265 1432 1267
rect 1426 1261 1428 1265
rect 1422 1259 1432 1261
rect 1426 1255 1428 1259
rect 1422 1253 1432 1255
rect 1426 1249 1428 1253
rect 1422 1247 1432 1249
rect 1426 1243 1428 1247
rect 1422 1181 1432 1243
rect 1426 1177 1428 1181
rect 1422 1175 1432 1177
rect 1426 1171 1428 1175
rect 1422 1169 1432 1171
rect 1426 1165 1428 1169
rect 1422 1163 1432 1165
rect 1426 1159 1428 1163
rect 1422 1157 1432 1159
rect 1426 1153 1428 1157
rect 96 1087 98 1091
rect 92 1085 102 1087
rect 96 1081 98 1085
rect 92 1079 102 1081
rect 96 1075 98 1079
rect 92 1073 102 1075
rect 96 1069 98 1073
rect 92 1067 102 1069
rect 96 1063 98 1067
rect 92 1001 102 1063
rect 96 997 98 1001
rect 92 995 102 997
rect 96 991 98 995
rect 92 989 102 991
rect 96 985 98 989
rect 92 983 102 985
rect 96 979 98 983
rect 92 977 102 979
rect 96 973 98 977
rect 92 911 102 973
rect 96 907 98 911
rect 92 905 102 907
rect 96 901 98 905
rect 92 899 102 901
rect 96 895 98 899
rect 92 893 102 895
rect 96 889 98 893
rect 92 887 102 889
rect 96 883 98 887
rect 92 821 102 883
rect 96 817 98 821
rect 92 815 102 817
rect 96 811 98 815
rect 92 809 102 811
rect 96 805 98 809
rect 92 803 102 805
rect 96 799 98 803
rect 92 797 102 799
rect 96 793 98 797
rect 92 731 102 793
rect 96 727 98 731
rect 92 725 102 727
rect 96 721 98 725
rect 92 719 102 721
rect 96 715 98 719
rect 92 713 102 715
rect 96 709 98 713
rect 92 707 102 709
rect 96 703 98 707
rect 92 641 102 703
rect 96 637 98 641
rect 92 635 102 637
rect 96 631 98 635
rect 92 629 102 631
rect 96 625 98 629
rect 92 623 102 625
rect 96 619 98 623
rect 92 617 102 619
rect 96 613 98 617
rect 92 551 102 613
rect 96 547 98 551
rect 92 545 102 547
rect 96 541 98 545
rect 92 539 102 541
rect 96 535 98 539
rect 92 533 102 535
rect 96 529 98 533
rect 92 527 102 529
rect 96 523 98 527
rect 92 461 102 523
rect 96 457 98 461
rect 92 455 102 457
rect 96 451 98 455
rect 92 449 102 451
rect 96 445 98 449
rect 92 443 102 445
rect 96 439 98 443
rect 92 437 102 439
rect 96 433 98 437
rect 92 371 102 433
rect 96 367 98 371
rect 92 365 102 367
rect 96 361 98 365
rect 92 359 102 361
rect 96 355 98 359
rect 92 353 102 355
rect 96 349 98 353
rect 92 347 102 349
rect 96 343 98 347
rect 92 281 102 343
rect 96 277 98 281
rect 92 275 102 277
rect 96 271 98 275
rect 92 269 102 271
rect 96 265 98 269
rect 92 263 102 265
rect 96 259 98 263
rect 92 257 102 259
rect 96 253 98 257
rect 92 191 102 253
rect 96 187 98 191
rect 92 185 102 187
rect 96 181 98 185
rect 92 179 102 181
rect 96 175 98 179
rect 92 173 102 175
rect 96 169 98 173
rect 92 167 102 169
rect 96 163 98 167
rect 92 126 102 163
rect 1422 1091 1432 1153
rect 1426 1087 1428 1091
rect 1422 1085 1432 1087
rect 1426 1081 1428 1085
rect 1422 1079 1432 1081
rect 1426 1075 1428 1079
rect 1422 1073 1432 1075
rect 1426 1069 1428 1073
rect 1422 1067 1432 1069
rect 1426 1063 1428 1067
rect 1422 1001 1432 1063
rect 1426 997 1428 1001
rect 1422 995 1432 997
rect 1426 991 1428 995
rect 1422 989 1432 991
rect 1426 985 1428 989
rect 1422 983 1432 985
rect 1426 979 1428 983
rect 1422 977 1432 979
rect 1426 973 1428 977
rect 1422 911 1432 973
rect 1426 907 1428 911
rect 1422 905 1432 907
rect 1426 901 1428 905
rect 1422 899 1432 901
rect 1426 895 1428 899
rect 1422 893 1432 895
rect 1426 889 1428 893
rect 1422 887 1432 889
rect 1426 883 1428 887
rect 1422 821 1432 883
rect 1426 817 1428 821
rect 1422 815 1432 817
rect 1426 811 1428 815
rect 1422 809 1432 811
rect 1426 805 1428 809
rect 1422 803 1432 805
rect 1426 799 1428 803
rect 1422 797 1432 799
rect 1426 793 1428 797
rect 1422 731 1432 793
rect 1426 727 1428 731
rect 1422 725 1432 727
rect 1426 721 1428 725
rect 1422 719 1432 721
rect 1426 715 1428 719
rect 1422 713 1432 715
rect 1426 709 1428 713
rect 1422 707 1432 709
rect 1426 703 1428 707
rect 1422 641 1432 703
rect 1426 637 1428 641
rect 1422 635 1432 637
rect 1426 631 1428 635
rect 1422 629 1432 631
rect 1426 625 1428 629
rect 1422 623 1432 625
rect 1426 619 1428 623
rect 1422 617 1432 619
rect 1426 613 1428 617
rect 1422 551 1432 613
rect 1426 547 1428 551
rect 1422 545 1432 547
rect 1426 541 1428 545
rect 1422 539 1432 541
rect 1426 535 1428 539
rect 1422 533 1432 535
rect 1426 529 1428 533
rect 1422 527 1432 529
rect 1426 523 1428 527
rect 1422 461 1432 523
rect 1426 457 1428 461
rect 1422 455 1432 457
rect 1426 451 1428 455
rect 1422 449 1432 451
rect 1426 445 1428 449
rect 1422 443 1432 445
rect 1426 439 1428 443
rect 1422 437 1432 439
rect 1426 433 1428 437
rect 1422 371 1432 433
rect 1426 367 1428 371
rect 1422 365 1432 367
rect 1426 361 1428 365
rect 1422 359 1432 361
rect 1426 355 1428 359
rect 1422 353 1432 355
rect 1426 349 1428 353
rect 1422 347 1432 349
rect 1426 343 1428 347
rect 1422 281 1432 343
rect 1426 277 1428 281
rect 1422 275 1432 277
rect 1426 271 1428 275
rect 1422 269 1432 271
rect 1426 265 1428 269
rect 1422 263 1432 265
rect 1426 259 1428 263
rect 1422 257 1432 259
rect 1426 253 1428 257
rect 1422 191 1432 253
rect 1426 187 1428 191
rect 1422 185 1432 187
rect 1426 181 1428 185
rect 1422 179 1432 181
rect 1426 175 1428 179
rect 1422 173 1432 175
rect 1426 169 1428 173
rect 1422 167 1432 169
rect 1426 163 1428 167
rect 1422 126 1432 163
rect 92 125 103 126
rect 1421 125 1432 126
rect 92 124 104 125
rect 1420 124 1432 125
rect 93 123 105 124
rect 1419 123 1431 124
rect 94 122 106 123
rect 1418 122 1430 123
rect 95 121 107 122
rect 1417 121 1429 122
rect 1438 121 1448 1403
rect 76 120 87 121
rect 96 120 108 121
rect 1416 120 1428 121
rect 1437 120 1448 121
rect 76 119 88 120
rect 97 119 109 120
rect 1415 119 1427 120
rect 1436 119 1448 120
rect 77 118 89 119
rect 98 118 110 119
rect 1414 118 1426 119
rect 1435 118 1447 119
rect 78 117 90 118
rect 99 117 111 118
rect 1413 117 1425 118
rect 1434 117 1446 118
rect 79 116 91 117
rect 100 116 112 117
rect 1412 116 1424 117
rect 1433 116 1445 117
rect 80 115 92 116
rect 101 115 113 116
rect 1411 115 1423 116
rect 1432 115 1444 116
rect 81 114 93 115
rect 102 114 114 115
rect 1410 114 1422 115
rect 1431 114 1443 115
rect 82 113 94 114
rect 103 113 115 114
rect 1409 113 1421 114
rect 1430 113 1442 114
rect 83 112 95 113
rect 104 112 116 113
rect 1408 112 1420 113
rect 1429 112 1441 113
rect 84 111 96 112
rect 105 111 117 112
rect 1407 111 1419 112
rect 1428 111 1440 112
rect 85 110 97 111
rect 106 110 118 111
rect 1406 110 1418 111
rect 1427 110 1439 111
rect 86 109 98 110
rect 107 109 119 110
rect 1405 109 1417 110
rect 1426 109 1438 110
rect 87 108 99 109
rect 108 108 120 109
rect 1404 108 1416 109
rect 1425 108 1437 109
rect 88 107 100 108
rect 109 107 121 108
rect 1403 107 1415 108
rect 1424 107 1436 108
rect 89 106 101 107
rect 110 106 122 107
rect 1402 106 1414 107
rect 1423 106 1435 107
rect 90 105 102 106
rect 111 105 123 106
rect 1401 105 1413 106
rect 1422 105 1434 106
rect 91 104 103 105
rect 112 104 124 105
rect 1400 104 1412 105
rect 1421 104 1433 105
rect 92 103 104 104
rect 113 103 125 104
rect 1399 103 1411 104
rect 1420 103 1432 104
rect 93 102 105 103
rect 114 102 126 103
rect 1398 102 1410 103
rect 1419 102 1431 103
rect 94 101 106 102
rect 115 101 163 102
rect 95 100 107 101
rect 116 100 163 101
rect 96 99 108 100
rect 117 99 163 100
rect 97 98 109 99
rect 118 98 163 99
rect 167 98 169 102
rect 173 98 175 102
rect 179 98 181 102
rect 185 98 187 102
rect 191 98 253 102
rect 257 98 259 102
rect 263 98 265 102
rect 269 98 271 102
rect 275 98 277 102
rect 281 98 343 102
rect 347 98 349 102
rect 353 98 355 102
rect 359 98 361 102
rect 365 98 367 102
rect 371 98 433 102
rect 437 98 439 102
rect 443 98 445 102
rect 449 98 451 102
rect 455 98 457 102
rect 461 98 523 102
rect 527 98 529 102
rect 533 98 535 102
rect 539 98 541 102
rect 545 98 547 102
rect 551 98 613 102
rect 617 98 619 102
rect 623 98 625 102
rect 629 98 631 102
rect 635 98 637 102
rect 641 98 703 102
rect 707 98 709 102
rect 713 98 715 102
rect 719 98 721 102
rect 725 98 727 102
rect 731 98 793 102
rect 797 98 799 102
rect 803 98 805 102
rect 809 98 811 102
rect 815 98 817 102
rect 821 98 883 102
rect 887 98 889 102
rect 893 98 895 102
rect 899 98 901 102
rect 905 98 907 102
rect 911 98 973 102
rect 977 98 979 102
rect 983 98 985 102
rect 989 98 991 102
rect 995 98 997 102
rect 1001 98 1063 102
rect 1067 98 1069 102
rect 1073 98 1075 102
rect 1079 98 1081 102
rect 1085 98 1087 102
rect 1091 98 1153 102
rect 1157 98 1159 102
rect 1163 98 1165 102
rect 1169 98 1171 102
rect 1175 98 1177 102
rect 1181 98 1243 102
rect 1247 98 1249 102
rect 1253 98 1255 102
rect 1259 98 1261 102
rect 1265 98 1267 102
rect 1271 98 1333 102
rect 1337 98 1339 102
rect 1343 98 1345 102
rect 1349 98 1351 102
rect 1355 98 1357 102
rect 1361 101 1409 102
rect 1418 101 1430 102
rect 1361 100 1408 101
rect 1417 100 1429 101
rect 1361 99 1407 100
rect 1416 99 1428 100
rect 1361 98 1406 99
rect 1415 98 1427 99
rect 98 97 110 98
rect 119 97 1405 98
rect 1414 97 1426 98
rect 99 96 111 97
rect 120 96 1404 97
rect 1413 96 1425 97
rect 100 95 112 96
rect 121 95 163 96
rect 101 94 113 95
rect 122 94 163 95
rect 102 93 114 94
rect 123 93 163 94
rect 103 92 115 93
rect 124 92 163 93
rect 167 92 169 96
rect 173 92 175 96
rect 179 92 181 96
rect 185 92 187 96
rect 191 92 253 96
rect 257 92 259 96
rect 263 92 265 96
rect 269 92 271 96
rect 275 92 277 96
rect 281 92 343 96
rect 347 92 349 96
rect 353 92 355 96
rect 359 92 361 96
rect 365 92 367 96
rect 371 92 433 96
rect 437 92 439 96
rect 443 92 445 96
rect 449 92 451 96
rect 455 92 457 96
rect 461 92 523 96
rect 527 92 529 96
rect 533 92 535 96
rect 539 92 541 96
rect 545 92 547 96
rect 551 92 613 96
rect 617 92 619 96
rect 623 92 625 96
rect 629 92 631 96
rect 635 92 637 96
rect 641 92 703 96
rect 707 92 709 96
rect 713 92 715 96
rect 719 92 721 96
rect 725 92 727 96
rect 731 92 793 96
rect 797 92 799 96
rect 803 92 805 96
rect 809 92 811 96
rect 815 92 817 96
rect 821 92 883 96
rect 887 92 889 96
rect 893 92 895 96
rect 899 92 901 96
rect 905 92 907 96
rect 911 92 973 96
rect 977 92 979 96
rect 983 92 985 96
rect 989 92 991 96
rect 995 92 997 96
rect 1001 92 1063 96
rect 1067 92 1069 96
rect 1073 92 1075 96
rect 1079 92 1081 96
rect 1085 92 1087 96
rect 1091 92 1153 96
rect 1157 92 1159 96
rect 1163 92 1165 96
rect 1169 92 1171 96
rect 1175 92 1177 96
rect 1181 92 1243 96
rect 1247 92 1249 96
rect 1253 92 1255 96
rect 1259 92 1261 96
rect 1265 92 1267 96
rect 1271 92 1333 96
rect 1337 92 1339 96
rect 1343 92 1345 96
rect 1349 92 1351 96
rect 1355 92 1357 96
rect 1361 95 1403 96
rect 1412 95 1424 96
rect 1361 94 1402 95
rect 1411 94 1423 95
rect 1361 93 1401 94
rect 1410 93 1422 94
rect 1361 92 1400 93
rect 1409 92 1421 93
rect 104 91 116 92
rect 1408 91 1420 92
rect 105 90 117 91
rect 1407 90 1419 91
rect 106 89 118 90
rect 1406 89 1418 90
rect 107 88 119 89
rect 1405 88 1417 89
rect 108 87 120 88
rect 1404 87 1416 88
rect 109 86 121 87
rect 1403 86 1415 87
rect 110 85 1414 86
rect 111 84 1413 85
rect 112 83 1412 84
rect 113 82 1411 83
rect 114 81 1410 82
rect 115 80 1409 81
rect 116 79 1408 80
rect 117 78 1407 79
rect 118 77 1406 78
rect 119 76 1405 77
<< metal2 >>
rect 162 1448 192 1454
rect 162 1444 163 1448
rect 167 1444 169 1448
rect 173 1444 175 1448
rect 179 1444 181 1448
rect 185 1444 187 1448
rect 191 1444 192 1448
rect 162 1442 192 1444
rect 162 1438 163 1442
rect 167 1438 169 1442
rect 173 1438 175 1442
rect 179 1438 181 1442
rect 185 1438 187 1442
rect 191 1438 192 1442
rect 162 1418 192 1438
rect 162 1414 163 1418
rect 167 1414 169 1418
rect 173 1414 175 1418
rect 179 1414 181 1418
rect 185 1414 187 1418
rect 191 1414 192 1418
rect 252 1414 282 1454
rect 342 1432 372 1454
rect 342 1428 343 1432
rect 347 1428 349 1432
rect 353 1428 355 1432
rect 359 1428 361 1432
rect 365 1428 367 1432
rect 371 1428 372 1432
rect 342 1426 372 1428
rect 342 1422 343 1426
rect 347 1422 349 1426
rect 353 1422 355 1426
rect 359 1422 361 1426
rect 365 1422 367 1426
rect 371 1422 372 1426
rect 342 1414 372 1422
rect 432 1432 462 1454
rect 432 1428 433 1432
rect 437 1428 439 1432
rect 443 1428 445 1432
rect 449 1428 451 1432
rect 455 1428 457 1432
rect 461 1428 462 1432
rect 432 1426 462 1428
rect 432 1422 433 1426
rect 437 1422 439 1426
rect 443 1422 445 1426
rect 449 1422 451 1426
rect 455 1422 457 1426
rect 461 1422 462 1426
rect 432 1414 462 1422
rect 522 1432 552 1454
rect 522 1428 523 1432
rect 527 1428 529 1432
rect 533 1428 535 1432
rect 539 1428 541 1432
rect 545 1428 547 1432
rect 551 1428 552 1432
rect 522 1426 552 1428
rect 522 1422 523 1426
rect 527 1422 529 1426
rect 533 1422 535 1426
rect 539 1422 541 1426
rect 545 1422 547 1426
rect 551 1422 552 1426
rect 522 1414 552 1422
rect 612 1432 642 1454
rect 612 1428 613 1432
rect 617 1428 619 1432
rect 623 1428 625 1432
rect 629 1428 631 1432
rect 635 1428 637 1432
rect 641 1428 642 1432
rect 612 1426 642 1428
rect 612 1422 613 1426
rect 617 1422 619 1426
rect 623 1422 625 1426
rect 629 1422 631 1426
rect 635 1422 637 1426
rect 641 1422 642 1426
rect 612 1414 642 1422
rect 702 1432 732 1454
rect 702 1428 703 1432
rect 707 1428 709 1432
rect 713 1428 715 1432
rect 719 1428 721 1432
rect 725 1428 727 1432
rect 731 1428 732 1432
rect 702 1426 732 1428
rect 702 1422 703 1426
rect 707 1422 709 1426
rect 713 1422 715 1426
rect 719 1422 721 1426
rect 725 1422 727 1426
rect 731 1422 732 1426
rect 702 1414 732 1422
rect 792 1432 822 1454
rect 792 1428 793 1432
rect 797 1428 799 1432
rect 803 1428 805 1432
rect 809 1428 811 1432
rect 815 1428 817 1432
rect 821 1428 822 1432
rect 792 1426 822 1428
rect 792 1422 793 1426
rect 797 1422 799 1426
rect 803 1422 805 1426
rect 809 1422 811 1426
rect 815 1422 817 1426
rect 821 1422 822 1426
rect 792 1414 822 1422
rect 882 1432 912 1454
rect 882 1428 883 1432
rect 887 1428 889 1432
rect 893 1428 895 1432
rect 899 1428 901 1432
rect 905 1428 907 1432
rect 911 1428 912 1432
rect 882 1426 912 1428
rect 882 1422 883 1426
rect 887 1422 889 1426
rect 893 1422 895 1426
rect 899 1422 901 1426
rect 905 1422 907 1426
rect 911 1422 912 1426
rect 882 1414 912 1422
rect 972 1432 1002 1454
rect 972 1428 973 1432
rect 977 1428 979 1432
rect 983 1428 985 1432
rect 989 1428 991 1432
rect 995 1428 997 1432
rect 1001 1428 1002 1432
rect 972 1426 1002 1428
rect 972 1422 973 1426
rect 977 1422 979 1426
rect 983 1422 985 1426
rect 989 1422 991 1426
rect 995 1422 997 1426
rect 1001 1422 1002 1426
rect 972 1414 1002 1422
rect 1062 1432 1092 1454
rect 1062 1428 1063 1432
rect 1067 1428 1069 1432
rect 1073 1428 1075 1432
rect 1079 1428 1081 1432
rect 1085 1428 1087 1432
rect 1091 1428 1092 1432
rect 1062 1426 1092 1428
rect 1062 1422 1063 1426
rect 1067 1422 1069 1426
rect 1073 1422 1075 1426
rect 1079 1422 1081 1426
rect 1085 1422 1087 1426
rect 1091 1422 1092 1426
rect 1062 1414 1092 1422
rect 1152 1432 1182 1454
rect 1152 1428 1153 1432
rect 1157 1428 1159 1432
rect 1163 1428 1165 1432
rect 1169 1428 1171 1432
rect 1175 1428 1177 1432
rect 1181 1428 1182 1432
rect 1152 1426 1182 1428
rect 1152 1422 1153 1426
rect 1157 1422 1159 1426
rect 1163 1422 1165 1426
rect 1169 1422 1171 1426
rect 1175 1422 1177 1426
rect 1181 1422 1182 1426
rect 1152 1414 1182 1422
rect 1242 1432 1272 1454
rect 1242 1428 1243 1432
rect 1247 1428 1249 1432
rect 1253 1428 1255 1432
rect 1259 1428 1261 1432
rect 1265 1428 1267 1432
rect 1271 1428 1272 1432
rect 1242 1426 1272 1428
rect 1242 1422 1243 1426
rect 1247 1422 1249 1426
rect 1253 1422 1255 1426
rect 1259 1422 1261 1426
rect 1265 1422 1267 1426
rect 1271 1422 1272 1426
rect 1242 1414 1272 1422
rect 1332 1432 1362 1454
rect 1332 1428 1333 1432
rect 1337 1428 1339 1432
rect 1343 1428 1345 1432
rect 1349 1428 1351 1432
rect 1355 1428 1357 1432
rect 1361 1428 1362 1432
rect 1332 1426 1362 1428
rect 1332 1422 1333 1426
rect 1337 1422 1339 1426
rect 1343 1422 1345 1426
rect 1349 1422 1351 1426
rect 1355 1422 1357 1426
rect 1361 1422 1362 1426
rect 1332 1414 1362 1422
rect 252 1407 271 1414
rect 187 1402 265 1407
rect 187 1383 192 1402
rect 174 1379 192 1383
rect 70 1360 114 1362
rect 70 1355 109 1360
rect 70 1352 114 1355
rect 70 1347 109 1352
rect 70 1344 114 1347
rect 70 1339 109 1344
rect 70 1332 114 1339
rect 1414 1361 1454 1362
rect 1414 1357 1422 1361
rect 1426 1357 1428 1361
rect 1432 1357 1454 1361
rect 1414 1355 1454 1357
rect 1414 1351 1422 1355
rect 1426 1351 1428 1355
rect 1432 1351 1454 1355
rect 1414 1349 1454 1351
rect 1414 1345 1422 1349
rect 1426 1345 1428 1349
rect 1432 1345 1454 1349
rect 1414 1343 1454 1345
rect 1414 1339 1422 1343
rect 1426 1339 1428 1343
rect 1432 1339 1454 1343
rect 1414 1337 1454 1339
rect 1414 1333 1422 1337
rect 1426 1333 1428 1337
rect 1432 1333 1454 1337
rect 1414 1332 1454 1333
rect 70 1271 115 1272
rect 70 1267 109 1271
rect 114 1267 115 1271
rect 70 1264 115 1267
rect 70 1260 109 1264
rect 114 1260 115 1264
rect 70 1257 115 1260
rect 70 1253 109 1257
rect 114 1253 115 1257
rect 70 1250 115 1253
rect 70 1246 109 1250
rect 114 1246 115 1250
rect 70 1242 115 1246
rect 1414 1271 1454 1272
rect 1414 1267 1422 1271
rect 1426 1267 1428 1271
rect 1432 1267 1454 1271
rect 1414 1265 1454 1267
rect 1414 1261 1422 1265
rect 1426 1261 1428 1265
rect 1432 1261 1454 1265
rect 1414 1259 1454 1261
rect 1414 1255 1422 1259
rect 1426 1255 1428 1259
rect 1432 1255 1454 1259
rect 1414 1253 1454 1255
rect 1414 1249 1422 1253
rect 1426 1249 1428 1253
rect 1432 1249 1454 1253
rect 1414 1247 1454 1249
rect 1414 1243 1422 1247
rect 1426 1243 1428 1247
rect 1432 1243 1454 1247
rect 1414 1242 1454 1243
rect 70 1178 124 1182
rect 70 1174 112 1178
rect 116 1174 119 1178
rect 123 1174 124 1178
rect 70 1171 124 1174
rect 70 1167 112 1171
rect 116 1167 119 1171
rect 123 1167 124 1171
rect 70 1165 124 1167
rect 70 1161 112 1165
rect 116 1161 119 1165
rect 123 1161 124 1165
rect 70 1159 124 1161
rect 70 1155 112 1159
rect 116 1155 119 1159
rect 123 1155 124 1159
rect 70 1152 124 1155
rect 1414 1181 1454 1182
rect 1414 1177 1422 1181
rect 1426 1177 1428 1181
rect 1432 1177 1454 1181
rect 1414 1175 1454 1177
rect 1414 1171 1422 1175
rect 1426 1171 1428 1175
rect 1432 1171 1454 1175
rect 1414 1169 1454 1171
rect 1414 1165 1422 1169
rect 1426 1165 1428 1169
rect 1432 1165 1454 1169
rect 1414 1163 1454 1165
rect 1414 1159 1422 1163
rect 1426 1159 1428 1163
rect 1432 1159 1454 1163
rect 1414 1157 1454 1159
rect 1414 1153 1422 1157
rect 1426 1153 1428 1157
rect 1432 1153 1454 1157
rect 1414 1152 1454 1153
rect 70 1091 110 1092
rect 70 1087 92 1091
rect 96 1087 98 1091
rect 102 1087 110 1091
rect 70 1085 110 1087
rect 70 1081 92 1085
rect 96 1081 98 1085
rect 102 1081 110 1085
rect 70 1079 110 1081
rect 70 1075 92 1079
rect 96 1075 98 1079
rect 102 1075 110 1079
rect 70 1073 110 1075
rect 70 1069 92 1073
rect 96 1069 98 1073
rect 102 1069 110 1073
rect 70 1067 110 1069
rect 70 1063 92 1067
rect 96 1063 98 1067
rect 102 1063 110 1067
rect 70 1062 110 1063
rect 1414 1091 1454 1092
rect 1414 1087 1422 1091
rect 1426 1087 1428 1091
rect 1432 1087 1454 1091
rect 1414 1085 1454 1087
rect 1414 1081 1422 1085
rect 1426 1081 1428 1085
rect 1432 1081 1454 1085
rect 1414 1079 1454 1081
rect 1414 1075 1422 1079
rect 1426 1075 1428 1079
rect 1432 1075 1454 1079
rect 1414 1073 1454 1075
rect 1414 1069 1422 1073
rect 1426 1069 1428 1073
rect 1432 1069 1454 1073
rect 1414 1067 1454 1069
rect 1414 1063 1422 1067
rect 1426 1063 1428 1067
rect 1432 1063 1454 1067
rect 1414 1062 1454 1063
rect 70 1001 110 1002
rect 70 997 92 1001
rect 96 997 98 1001
rect 102 997 110 1001
rect 70 995 110 997
rect 70 991 92 995
rect 96 991 98 995
rect 102 991 110 995
rect 70 989 110 991
rect 70 985 92 989
rect 96 985 98 989
rect 102 985 110 989
rect 70 983 110 985
rect 70 979 92 983
rect 96 979 98 983
rect 102 979 110 983
rect 70 977 110 979
rect 70 973 92 977
rect 96 973 98 977
rect 102 973 110 977
rect 70 972 110 973
rect 1414 1001 1454 1002
rect 1414 997 1422 1001
rect 1426 997 1428 1001
rect 1432 997 1454 1001
rect 1414 995 1454 997
rect 1414 991 1422 995
rect 1426 991 1428 995
rect 1432 991 1454 995
rect 1414 989 1454 991
rect 1414 985 1422 989
rect 1426 985 1428 989
rect 1432 985 1454 989
rect 1414 983 1454 985
rect 1414 979 1422 983
rect 1426 979 1428 983
rect 1432 979 1454 983
rect 1414 977 1454 979
rect 1414 973 1422 977
rect 1426 973 1428 977
rect 1432 973 1454 977
rect 1414 972 1454 973
rect 70 911 110 912
rect 70 907 92 911
rect 96 907 98 911
rect 102 907 110 911
rect 70 905 110 907
rect 70 901 92 905
rect 96 901 98 905
rect 102 901 110 905
rect 70 899 110 901
rect 70 895 92 899
rect 96 895 98 899
rect 102 895 110 899
rect 70 893 110 895
rect 70 889 92 893
rect 96 889 98 893
rect 102 889 110 893
rect 70 887 110 889
rect 70 883 92 887
rect 96 883 98 887
rect 102 883 110 887
rect 70 882 110 883
rect 1414 911 1454 912
rect 1414 907 1422 911
rect 1426 907 1428 911
rect 1432 907 1454 911
rect 1414 905 1454 907
rect 1414 901 1422 905
rect 1426 901 1428 905
rect 1432 901 1454 905
rect 1414 899 1454 901
rect 1414 895 1422 899
rect 1426 895 1428 899
rect 1432 895 1454 899
rect 1414 893 1454 895
rect 1414 889 1422 893
rect 1426 889 1428 893
rect 1432 889 1454 893
rect 1414 887 1454 889
rect 1414 883 1422 887
rect 1426 883 1428 887
rect 1432 883 1454 887
rect 1414 882 1454 883
rect 70 821 110 822
rect 70 817 92 821
rect 96 817 98 821
rect 102 817 110 821
rect 70 815 110 817
rect 70 811 92 815
rect 96 811 98 815
rect 102 811 110 815
rect 70 809 110 811
rect 70 805 92 809
rect 96 805 98 809
rect 102 805 110 809
rect 70 803 110 805
rect 70 799 92 803
rect 96 799 98 803
rect 102 799 110 803
rect 70 797 110 799
rect 70 793 92 797
rect 96 793 98 797
rect 102 793 110 797
rect 70 792 110 793
rect 1414 821 1454 822
rect 1414 817 1422 821
rect 1426 817 1428 821
rect 1432 817 1454 821
rect 1414 815 1454 817
rect 1414 811 1422 815
rect 1426 811 1428 815
rect 1432 811 1454 815
rect 1414 809 1454 811
rect 1414 805 1422 809
rect 1426 805 1428 809
rect 1432 805 1454 809
rect 1414 803 1454 805
rect 1414 799 1422 803
rect 1426 799 1428 803
rect 1432 799 1454 803
rect 1414 797 1454 799
rect 1414 793 1422 797
rect 1426 793 1428 797
rect 1432 793 1454 797
rect 1414 792 1454 793
rect 70 731 110 732
rect 70 727 92 731
rect 96 727 98 731
rect 102 727 110 731
rect 70 725 110 727
rect 70 721 92 725
rect 96 721 98 725
rect 102 721 110 725
rect 70 719 110 721
rect 70 715 92 719
rect 96 715 98 719
rect 102 715 110 719
rect 70 713 110 715
rect 70 709 92 713
rect 96 709 98 713
rect 102 709 110 713
rect 70 707 110 709
rect 70 703 92 707
rect 96 703 98 707
rect 102 703 110 707
rect 70 702 110 703
rect 1414 731 1454 732
rect 1414 727 1422 731
rect 1426 727 1428 731
rect 1432 727 1454 731
rect 1414 725 1454 727
rect 1414 721 1422 725
rect 1426 721 1428 725
rect 1432 721 1454 725
rect 1414 719 1454 721
rect 1414 715 1422 719
rect 1426 715 1428 719
rect 1432 715 1454 719
rect 1414 713 1454 715
rect 1414 709 1422 713
rect 1426 709 1428 713
rect 1432 709 1454 713
rect 1414 707 1454 709
rect 1414 703 1422 707
rect 1426 703 1428 707
rect 1432 703 1454 707
rect 1414 702 1454 703
rect 70 641 110 642
rect 70 637 92 641
rect 96 637 98 641
rect 102 637 110 641
rect 70 635 110 637
rect 70 631 92 635
rect 96 631 98 635
rect 102 631 110 635
rect 70 629 110 631
rect 70 625 92 629
rect 96 625 98 629
rect 102 625 110 629
rect 70 623 110 625
rect 70 619 92 623
rect 96 619 98 623
rect 102 619 110 623
rect 70 617 110 619
rect 70 613 92 617
rect 96 613 98 617
rect 102 613 110 617
rect 70 612 110 613
rect 1414 641 1454 642
rect 1414 637 1422 641
rect 1426 637 1428 641
rect 1432 637 1454 641
rect 1414 635 1454 637
rect 1414 631 1422 635
rect 1426 631 1428 635
rect 1432 631 1454 635
rect 1414 629 1454 631
rect 1414 625 1422 629
rect 1426 625 1428 629
rect 1432 625 1454 629
rect 1414 623 1454 625
rect 1414 619 1422 623
rect 1426 619 1428 623
rect 1432 619 1454 623
rect 1414 617 1454 619
rect 1414 613 1422 617
rect 1426 613 1428 617
rect 1432 613 1454 617
rect 1414 612 1454 613
rect 70 551 110 552
rect 70 547 92 551
rect 96 547 98 551
rect 102 547 110 551
rect 70 545 110 547
rect 70 541 92 545
rect 96 541 98 545
rect 102 541 110 545
rect 70 539 110 541
rect 70 535 92 539
rect 96 535 98 539
rect 102 535 110 539
rect 70 533 110 535
rect 70 529 92 533
rect 96 529 98 533
rect 102 529 110 533
rect 70 527 110 529
rect 70 523 92 527
rect 96 523 98 527
rect 102 523 110 527
rect 70 522 110 523
rect 1414 551 1454 552
rect 1414 547 1422 551
rect 1426 547 1428 551
rect 1432 547 1454 551
rect 1414 545 1454 547
rect 1414 541 1422 545
rect 1426 541 1428 545
rect 1432 541 1454 545
rect 1414 539 1454 541
rect 1414 535 1422 539
rect 1426 535 1428 539
rect 1432 535 1454 539
rect 1414 533 1454 535
rect 1414 529 1422 533
rect 1426 529 1428 533
rect 1432 529 1454 533
rect 1414 527 1454 529
rect 1414 523 1422 527
rect 1426 523 1428 527
rect 1432 523 1454 527
rect 1414 522 1454 523
rect 70 461 110 462
rect 70 457 92 461
rect 96 457 98 461
rect 102 457 110 461
rect 70 455 110 457
rect 70 451 92 455
rect 96 451 98 455
rect 102 451 110 455
rect 70 449 110 451
rect 70 445 92 449
rect 96 445 98 449
rect 102 445 110 449
rect 70 443 110 445
rect 70 439 92 443
rect 96 439 98 443
rect 102 439 110 443
rect 70 437 110 439
rect 70 433 92 437
rect 96 433 98 437
rect 102 433 110 437
rect 70 432 110 433
rect 1414 461 1454 462
rect 1414 457 1422 461
rect 1426 457 1428 461
rect 1432 457 1454 461
rect 1414 455 1454 457
rect 1414 451 1422 455
rect 1426 451 1428 455
rect 1432 451 1454 455
rect 1414 449 1454 451
rect 1414 445 1422 449
rect 1426 445 1428 449
rect 1432 445 1454 449
rect 1414 443 1454 445
rect 1414 439 1422 443
rect 1426 439 1428 443
rect 1432 439 1454 443
rect 1414 437 1454 439
rect 1414 433 1422 437
rect 1426 433 1428 437
rect 1432 433 1454 437
rect 1414 432 1454 433
rect 70 371 110 372
rect 70 367 92 371
rect 96 367 98 371
rect 102 367 110 371
rect 70 365 110 367
rect 70 361 92 365
rect 96 361 98 365
rect 102 361 110 365
rect 70 359 110 361
rect 70 355 92 359
rect 96 355 98 359
rect 102 355 110 359
rect 70 353 110 355
rect 70 349 92 353
rect 96 349 98 353
rect 102 349 110 353
rect 70 347 110 349
rect 70 343 92 347
rect 96 343 98 347
rect 102 343 110 347
rect 70 342 110 343
rect 1414 371 1454 372
rect 1414 367 1422 371
rect 1426 367 1428 371
rect 1432 367 1454 371
rect 1414 365 1454 367
rect 1414 361 1422 365
rect 1426 361 1428 365
rect 1432 361 1454 365
rect 1414 359 1454 361
rect 1414 355 1422 359
rect 1426 355 1428 359
rect 1432 355 1454 359
rect 1414 353 1454 355
rect 1414 349 1422 353
rect 1426 349 1428 353
rect 1432 349 1454 353
rect 1414 347 1454 349
rect 1414 343 1422 347
rect 1426 343 1428 347
rect 1432 343 1454 347
rect 1414 342 1454 343
rect 70 281 110 282
rect 70 277 92 281
rect 96 277 98 281
rect 102 277 110 281
rect 70 275 110 277
rect 70 271 92 275
rect 96 271 98 275
rect 102 271 110 275
rect 70 269 110 271
rect 70 265 92 269
rect 96 265 98 269
rect 102 265 110 269
rect 70 263 110 265
rect 70 259 92 263
rect 96 259 98 263
rect 102 259 110 263
rect 70 257 110 259
rect 70 253 92 257
rect 96 253 98 257
rect 102 253 110 257
rect 70 252 110 253
rect 1414 281 1454 282
rect 1414 277 1422 281
rect 1426 277 1428 281
rect 1432 277 1454 281
rect 1414 275 1454 277
rect 1414 271 1422 275
rect 1426 271 1428 275
rect 1432 271 1454 275
rect 1414 269 1454 271
rect 1414 265 1422 269
rect 1426 265 1428 269
rect 1432 265 1454 269
rect 1414 263 1454 265
rect 1414 259 1422 263
rect 1426 259 1428 263
rect 1432 259 1454 263
rect 1414 257 1454 259
rect 1414 253 1422 257
rect 1426 253 1428 257
rect 1432 253 1454 257
rect 1414 252 1454 253
rect 70 191 110 192
rect 70 187 92 191
rect 96 187 98 191
rect 102 187 110 191
rect 70 185 110 187
rect 70 181 92 185
rect 96 181 98 185
rect 102 181 110 185
rect 70 179 110 181
rect 70 175 92 179
rect 96 175 98 179
rect 102 175 110 179
rect 70 173 110 175
rect 70 169 92 173
rect 96 169 98 173
rect 102 169 110 173
rect 70 167 110 169
rect 70 163 92 167
rect 96 163 98 167
rect 102 163 110 167
rect 70 162 110 163
rect 1414 191 1454 192
rect 1414 187 1422 191
rect 1426 187 1428 191
rect 1432 187 1454 191
rect 1414 185 1454 187
rect 1414 181 1422 185
rect 1426 181 1428 185
rect 1432 181 1454 185
rect 1414 179 1454 181
rect 1414 175 1422 179
rect 1426 175 1428 179
rect 1432 175 1454 179
rect 1414 173 1454 175
rect 1414 169 1422 173
rect 1426 169 1428 173
rect 1432 169 1454 173
rect 1414 167 1454 169
rect 1414 163 1422 167
rect 1426 163 1428 167
rect 1432 163 1454 167
rect 1414 162 1454 163
rect 162 102 192 110
rect 162 98 163 102
rect 167 98 169 102
rect 173 98 175 102
rect 179 98 181 102
rect 185 98 187 102
rect 191 98 192 102
rect 162 96 192 98
rect 162 92 163 96
rect 167 92 169 96
rect 173 92 175 96
rect 179 92 181 96
rect 185 92 187 96
rect 191 92 192 96
rect 162 70 192 92
rect 252 102 282 110
rect 252 98 253 102
rect 257 98 259 102
rect 263 98 265 102
rect 269 98 271 102
rect 275 98 277 102
rect 281 98 282 102
rect 252 96 282 98
rect 252 92 253 96
rect 257 92 259 96
rect 263 92 265 96
rect 269 92 271 96
rect 275 92 277 96
rect 281 92 282 96
rect 252 70 282 92
rect 342 102 372 110
rect 342 98 343 102
rect 347 98 349 102
rect 353 98 355 102
rect 359 98 361 102
rect 365 98 367 102
rect 371 98 372 102
rect 342 96 372 98
rect 342 92 343 96
rect 347 92 349 96
rect 353 92 355 96
rect 359 92 361 96
rect 365 92 367 96
rect 371 92 372 96
rect 342 70 372 92
rect 432 102 462 110
rect 432 98 433 102
rect 437 98 439 102
rect 443 98 445 102
rect 449 98 451 102
rect 455 98 457 102
rect 461 98 462 102
rect 432 96 462 98
rect 432 92 433 96
rect 437 92 439 96
rect 443 92 445 96
rect 449 92 451 96
rect 455 92 457 96
rect 461 92 462 96
rect 432 70 462 92
rect 522 102 552 110
rect 522 98 523 102
rect 527 98 529 102
rect 533 98 535 102
rect 539 98 541 102
rect 545 98 547 102
rect 551 98 552 102
rect 522 96 552 98
rect 522 92 523 96
rect 527 92 529 96
rect 533 92 535 96
rect 539 92 541 96
rect 545 92 547 96
rect 551 92 552 96
rect 522 70 552 92
rect 612 102 642 110
rect 612 98 613 102
rect 617 98 619 102
rect 623 98 625 102
rect 629 98 631 102
rect 635 98 637 102
rect 641 98 642 102
rect 612 96 642 98
rect 612 92 613 96
rect 617 92 619 96
rect 623 92 625 96
rect 629 92 631 96
rect 635 92 637 96
rect 641 92 642 96
rect 612 70 642 92
rect 702 102 732 110
rect 702 98 703 102
rect 707 98 709 102
rect 713 98 715 102
rect 719 98 721 102
rect 725 98 727 102
rect 731 98 732 102
rect 702 96 732 98
rect 702 92 703 96
rect 707 92 709 96
rect 713 92 715 96
rect 719 92 721 96
rect 725 92 727 96
rect 731 92 732 96
rect 702 70 732 92
rect 792 102 822 110
rect 792 98 793 102
rect 797 98 799 102
rect 803 98 805 102
rect 809 98 811 102
rect 815 98 817 102
rect 821 98 822 102
rect 792 96 822 98
rect 792 92 793 96
rect 797 92 799 96
rect 803 92 805 96
rect 809 92 811 96
rect 815 92 817 96
rect 821 92 822 96
rect 792 70 822 92
rect 882 102 912 110
rect 882 98 883 102
rect 887 98 889 102
rect 893 98 895 102
rect 899 98 901 102
rect 905 98 907 102
rect 911 98 912 102
rect 882 96 912 98
rect 882 92 883 96
rect 887 92 889 96
rect 893 92 895 96
rect 899 92 901 96
rect 905 92 907 96
rect 911 92 912 96
rect 882 70 912 92
rect 972 102 1002 110
rect 972 98 973 102
rect 977 98 979 102
rect 983 98 985 102
rect 989 98 991 102
rect 995 98 997 102
rect 1001 98 1002 102
rect 972 96 1002 98
rect 972 92 973 96
rect 977 92 979 96
rect 983 92 985 96
rect 989 92 991 96
rect 995 92 997 96
rect 1001 92 1002 96
rect 972 70 1002 92
rect 1062 102 1092 110
rect 1062 98 1063 102
rect 1067 98 1069 102
rect 1073 98 1075 102
rect 1079 98 1081 102
rect 1085 98 1087 102
rect 1091 98 1092 102
rect 1062 96 1092 98
rect 1062 92 1063 96
rect 1067 92 1069 96
rect 1073 92 1075 96
rect 1079 92 1081 96
rect 1085 92 1087 96
rect 1091 92 1092 96
rect 1062 70 1092 92
rect 1152 102 1182 110
rect 1152 98 1153 102
rect 1157 98 1159 102
rect 1163 98 1165 102
rect 1169 98 1171 102
rect 1175 98 1177 102
rect 1181 98 1182 102
rect 1152 96 1182 98
rect 1152 92 1153 96
rect 1157 92 1159 96
rect 1163 92 1165 96
rect 1169 92 1171 96
rect 1175 92 1177 96
rect 1181 92 1182 96
rect 1152 70 1182 92
rect 1242 102 1272 110
rect 1242 98 1243 102
rect 1247 98 1249 102
rect 1253 98 1255 102
rect 1259 98 1261 102
rect 1265 98 1267 102
rect 1271 98 1272 102
rect 1242 96 1272 98
rect 1242 92 1243 96
rect 1247 92 1249 96
rect 1253 92 1255 96
rect 1259 92 1261 96
rect 1265 92 1267 96
rect 1271 92 1272 96
rect 1242 70 1272 92
rect 1332 102 1362 110
rect 1332 98 1333 102
rect 1337 98 1339 102
rect 1343 98 1345 102
rect 1349 98 1351 102
rect 1355 98 1357 102
rect 1361 98 1362 102
rect 1332 96 1362 98
rect 1332 92 1333 96
rect 1337 92 1339 96
rect 1343 92 1345 96
rect 1349 92 1351 96
rect 1355 92 1357 96
rect 1361 92 1362 96
rect 1332 70 1362 92
<< polycontact >>
rect 135 1391 139 1395
rect 116 1339 120 1359
rect 154 1353 158 1357
rect 162 1353 166 1357
<< m2contact >>
rect 163 1444 167 1448
rect 169 1444 173 1448
rect 175 1444 179 1448
rect 181 1444 185 1448
rect 187 1444 191 1448
rect 163 1438 167 1442
rect 169 1438 173 1442
rect 175 1438 179 1442
rect 181 1438 185 1442
rect 187 1438 191 1442
rect 343 1428 347 1432
rect 349 1428 353 1432
rect 355 1428 359 1432
rect 361 1428 365 1432
rect 367 1428 371 1432
rect 433 1428 437 1432
rect 439 1428 443 1432
rect 445 1428 449 1432
rect 451 1428 455 1432
rect 457 1428 461 1432
rect 523 1428 527 1432
rect 529 1428 533 1432
rect 535 1428 539 1432
rect 541 1428 545 1432
rect 547 1428 551 1432
rect 613 1428 617 1432
rect 619 1428 623 1432
rect 625 1428 629 1432
rect 631 1428 635 1432
rect 637 1428 641 1432
rect 703 1428 707 1432
rect 709 1428 713 1432
rect 715 1428 719 1432
rect 721 1428 725 1432
rect 727 1428 731 1432
rect 793 1428 797 1432
rect 799 1428 803 1432
rect 805 1428 809 1432
rect 811 1428 815 1432
rect 817 1428 821 1432
rect 883 1428 887 1432
rect 889 1428 893 1432
rect 895 1428 899 1432
rect 901 1428 905 1432
rect 907 1428 911 1432
rect 973 1428 977 1432
rect 979 1428 983 1432
rect 985 1428 989 1432
rect 991 1428 995 1432
rect 997 1428 1001 1432
rect 1063 1428 1067 1432
rect 1069 1428 1073 1432
rect 1075 1428 1079 1432
rect 1081 1428 1085 1432
rect 1087 1428 1091 1432
rect 1153 1428 1157 1432
rect 1159 1428 1163 1432
rect 1165 1428 1169 1432
rect 1171 1428 1175 1432
rect 1177 1428 1181 1432
rect 1243 1428 1247 1432
rect 1249 1428 1253 1432
rect 1255 1428 1259 1432
rect 1261 1428 1265 1432
rect 1267 1428 1271 1432
rect 1333 1428 1337 1432
rect 1339 1428 1343 1432
rect 1345 1428 1349 1432
rect 1351 1428 1355 1432
rect 1357 1428 1361 1432
rect 343 1422 347 1426
rect 349 1422 353 1426
rect 355 1422 359 1426
rect 361 1422 365 1426
rect 367 1422 371 1426
rect 433 1422 437 1426
rect 439 1422 443 1426
rect 445 1422 449 1426
rect 451 1422 455 1426
rect 457 1422 461 1426
rect 523 1422 527 1426
rect 529 1422 533 1426
rect 535 1422 539 1426
rect 541 1422 545 1426
rect 547 1422 551 1426
rect 613 1422 617 1426
rect 619 1422 623 1426
rect 625 1422 629 1426
rect 631 1422 635 1426
rect 637 1422 641 1426
rect 703 1422 707 1426
rect 709 1422 713 1426
rect 715 1422 719 1426
rect 721 1422 725 1426
rect 727 1422 731 1426
rect 793 1422 797 1426
rect 799 1422 803 1426
rect 805 1422 809 1426
rect 811 1422 815 1426
rect 817 1422 821 1426
rect 883 1422 887 1426
rect 889 1422 893 1426
rect 895 1422 899 1426
rect 901 1422 905 1426
rect 907 1422 911 1426
rect 973 1422 977 1426
rect 979 1422 983 1426
rect 985 1422 989 1426
rect 991 1422 995 1426
rect 997 1422 1001 1426
rect 1063 1422 1067 1426
rect 1069 1422 1073 1426
rect 1075 1422 1079 1426
rect 1081 1422 1085 1426
rect 1087 1422 1091 1426
rect 1153 1422 1157 1426
rect 1159 1422 1163 1426
rect 1165 1422 1169 1426
rect 1171 1422 1175 1426
rect 1177 1422 1181 1426
rect 1243 1422 1247 1426
rect 1249 1422 1253 1426
rect 1255 1422 1259 1426
rect 1261 1422 1265 1426
rect 1267 1422 1271 1426
rect 1333 1422 1337 1426
rect 1339 1422 1343 1426
rect 1345 1422 1349 1426
rect 1351 1422 1355 1426
rect 1357 1422 1361 1426
rect 163 1414 167 1418
rect 169 1414 173 1418
rect 175 1414 179 1418
rect 181 1414 185 1418
rect 187 1414 191 1418
rect 170 1379 174 1383
rect 109 1355 114 1360
rect 109 1347 114 1352
rect 109 1339 114 1344
rect 1422 1357 1426 1361
rect 1428 1357 1432 1361
rect 1422 1351 1426 1355
rect 1428 1351 1432 1355
rect 1422 1345 1426 1349
rect 1428 1345 1432 1349
rect 1422 1339 1426 1343
rect 1428 1339 1432 1343
rect 109 1267 114 1271
rect 109 1260 114 1264
rect 109 1253 114 1257
rect 109 1246 114 1250
rect 1422 1333 1426 1337
rect 1428 1333 1432 1337
rect 112 1174 116 1178
rect 119 1174 123 1178
rect 112 1167 116 1171
rect 119 1167 123 1171
rect 112 1161 116 1165
rect 119 1161 123 1165
rect 112 1155 116 1159
rect 119 1155 123 1159
rect 1422 1267 1426 1271
rect 1428 1267 1432 1271
rect 1422 1261 1426 1265
rect 1428 1261 1432 1265
rect 1422 1255 1426 1259
rect 1428 1255 1432 1259
rect 1422 1249 1426 1253
rect 1428 1249 1432 1253
rect 1422 1243 1426 1247
rect 1428 1243 1432 1247
rect 1422 1177 1426 1181
rect 1428 1177 1432 1181
rect 1422 1171 1426 1175
rect 1428 1171 1432 1175
rect 1422 1165 1426 1169
rect 1428 1165 1432 1169
rect 1422 1159 1426 1163
rect 1428 1159 1432 1163
rect 1422 1153 1426 1157
rect 1428 1153 1432 1157
rect 92 1087 96 1091
rect 98 1087 102 1091
rect 92 1081 96 1085
rect 98 1081 102 1085
rect 92 1075 96 1079
rect 98 1075 102 1079
rect 92 1069 96 1073
rect 98 1069 102 1073
rect 92 1063 96 1067
rect 98 1063 102 1067
rect 92 997 96 1001
rect 98 997 102 1001
rect 92 991 96 995
rect 98 991 102 995
rect 92 985 96 989
rect 98 985 102 989
rect 92 979 96 983
rect 98 979 102 983
rect 92 973 96 977
rect 98 973 102 977
rect 92 907 96 911
rect 98 907 102 911
rect 92 901 96 905
rect 98 901 102 905
rect 92 895 96 899
rect 98 895 102 899
rect 92 889 96 893
rect 98 889 102 893
rect 92 883 96 887
rect 98 883 102 887
rect 92 817 96 821
rect 98 817 102 821
rect 92 811 96 815
rect 98 811 102 815
rect 92 805 96 809
rect 98 805 102 809
rect 92 799 96 803
rect 98 799 102 803
rect 92 793 96 797
rect 98 793 102 797
rect 92 727 96 731
rect 98 727 102 731
rect 92 721 96 725
rect 98 721 102 725
rect 92 715 96 719
rect 98 715 102 719
rect 92 709 96 713
rect 98 709 102 713
rect 92 703 96 707
rect 98 703 102 707
rect 92 637 96 641
rect 98 637 102 641
rect 92 631 96 635
rect 98 631 102 635
rect 92 625 96 629
rect 98 625 102 629
rect 92 619 96 623
rect 98 619 102 623
rect 92 613 96 617
rect 98 613 102 617
rect 92 547 96 551
rect 98 547 102 551
rect 92 541 96 545
rect 98 541 102 545
rect 92 535 96 539
rect 98 535 102 539
rect 92 529 96 533
rect 98 529 102 533
rect 92 523 96 527
rect 98 523 102 527
rect 92 457 96 461
rect 98 457 102 461
rect 92 451 96 455
rect 98 451 102 455
rect 92 445 96 449
rect 98 445 102 449
rect 92 439 96 443
rect 98 439 102 443
rect 92 433 96 437
rect 98 433 102 437
rect 92 367 96 371
rect 98 367 102 371
rect 92 361 96 365
rect 98 361 102 365
rect 92 355 96 359
rect 98 355 102 359
rect 92 349 96 353
rect 98 349 102 353
rect 92 343 96 347
rect 98 343 102 347
rect 92 277 96 281
rect 98 277 102 281
rect 92 271 96 275
rect 98 271 102 275
rect 92 265 96 269
rect 98 265 102 269
rect 92 259 96 263
rect 98 259 102 263
rect 92 253 96 257
rect 98 253 102 257
rect 92 187 96 191
rect 98 187 102 191
rect 92 181 96 185
rect 98 181 102 185
rect 92 175 96 179
rect 98 175 102 179
rect 92 169 96 173
rect 98 169 102 173
rect 92 163 96 167
rect 98 163 102 167
rect 1422 1087 1426 1091
rect 1428 1087 1432 1091
rect 1422 1081 1426 1085
rect 1428 1081 1432 1085
rect 1422 1075 1426 1079
rect 1428 1075 1432 1079
rect 1422 1069 1426 1073
rect 1428 1069 1432 1073
rect 1422 1063 1426 1067
rect 1428 1063 1432 1067
rect 1422 997 1426 1001
rect 1428 997 1432 1001
rect 1422 991 1426 995
rect 1428 991 1432 995
rect 1422 985 1426 989
rect 1428 985 1432 989
rect 1422 979 1426 983
rect 1428 979 1432 983
rect 1422 973 1426 977
rect 1428 973 1432 977
rect 1422 907 1426 911
rect 1428 907 1432 911
rect 1422 901 1426 905
rect 1428 901 1432 905
rect 1422 895 1426 899
rect 1428 895 1432 899
rect 1422 889 1426 893
rect 1428 889 1432 893
rect 1422 883 1426 887
rect 1428 883 1432 887
rect 1422 817 1426 821
rect 1428 817 1432 821
rect 1422 811 1426 815
rect 1428 811 1432 815
rect 1422 805 1426 809
rect 1428 805 1432 809
rect 1422 799 1426 803
rect 1428 799 1432 803
rect 1422 793 1426 797
rect 1428 793 1432 797
rect 1422 727 1426 731
rect 1428 727 1432 731
rect 1422 721 1426 725
rect 1428 721 1432 725
rect 1422 715 1426 719
rect 1428 715 1432 719
rect 1422 709 1426 713
rect 1428 709 1432 713
rect 1422 703 1426 707
rect 1428 703 1432 707
rect 1422 637 1426 641
rect 1428 637 1432 641
rect 1422 631 1426 635
rect 1428 631 1432 635
rect 1422 625 1426 629
rect 1428 625 1432 629
rect 1422 619 1426 623
rect 1428 619 1432 623
rect 1422 613 1426 617
rect 1428 613 1432 617
rect 1422 547 1426 551
rect 1428 547 1432 551
rect 1422 541 1426 545
rect 1428 541 1432 545
rect 1422 535 1426 539
rect 1428 535 1432 539
rect 1422 529 1426 533
rect 1428 529 1432 533
rect 1422 523 1426 527
rect 1428 523 1432 527
rect 1422 457 1426 461
rect 1428 457 1432 461
rect 1422 451 1426 455
rect 1428 451 1432 455
rect 1422 445 1426 449
rect 1428 445 1432 449
rect 1422 439 1426 443
rect 1428 439 1432 443
rect 1422 433 1426 437
rect 1428 433 1432 437
rect 1422 367 1426 371
rect 1428 367 1432 371
rect 1422 361 1426 365
rect 1428 361 1432 365
rect 1422 355 1426 359
rect 1428 355 1432 359
rect 1422 349 1426 353
rect 1428 349 1432 353
rect 1422 343 1426 347
rect 1428 343 1432 347
rect 1422 277 1426 281
rect 1428 277 1432 281
rect 1422 271 1426 275
rect 1428 271 1432 275
rect 1422 265 1426 269
rect 1428 265 1432 269
rect 1422 259 1426 263
rect 1428 259 1432 263
rect 1422 253 1426 257
rect 1428 253 1432 257
rect 1422 187 1426 191
rect 1428 187 1432 191
rect 1422 181 1426 185
rect 1428 181 1432 185
rect 1422 175 1426 179
rect 1428 175 1432 179
rect 1422 169 1426 173
rect 1428 169 1432 173
rect 1422 163 1426 167
rect 1428 163 1432 167
rect 163 98 167 102
rect 169 98 173 102
rect 175 98 179 102
rect 181 98 185 102
rect 187 98 191 102
rect 253 98 257 102
rect 259 98 263 102
rect 265 98 269 102
rect 271 98 275 102
rect 277 98 281 102
rect 343 98 347 102
rect 349 98 353 102
rect 355 98 359 102
rect 361 98 365 102
rect 367 98 371 102
rect 433 98 437 102
rect 439 98 443 102
rect 445 98 449 102
rect 451 98 455 102
rect 457 98 461 102
rect 523 98 527 102
rect 529 98 533 102
rect 535 98 539 102
rect 541 98 545 102
rect 547 98 551 102
rect 613 98 617 102
rect 619 98 623 102
rect 625 98 629 102
rect 631 98 635 102
rect 637 98 641 102
rect 703 98 707 102
rect 709 98 713 102
rect 715 98 719 102
rect 721 98 725 102
rect 727 98 731 102
rect 793 98 797 102
rect 799 98 803 102
rect 805 98 809 102
rect 811 98 815 102
rect 817 98 821 102
rect 883 98 887 102
rect 889 98 893 102
rect 895 98 899 102
rect 901 98 905 102
rect 907 98 911 102
rect 973 98 977 102
rect 979 98 983 102
rect 985 98 989 102
rect 991 98 995 102
rect 997 98 1001 102
rect 1063 98 1067 102
rect 1069 98 1073 102
rect 1075 98 1079 102
rect 1081 98 1085 102
rect 1087 98 1091 102
rect 1153 98 1157 102
rect 1159 98 1163 102
rect 1165 98 1169 102
rect 1171 98 1175 102
rect 1177 98 1181 102
rect 1243 98 1247 102
rect 1249 98 1253 102
rect 1255 98 1259 102
rect 1261 98 1265 102
rect 1267 98 1271 102
rect 1333 98 1337 102
rect 1339 98 1343 102
rect 1345 98 1349 102
rect 1351 98 1355 102
rect 1357 98 1361 102
rect 163 92 167 96
rect 169 92 173 96
rect 175 92 179 96
rect 181 92 185 96
rect 187 92 191 96
rect 253 92 257 96
rect 259 92 263 96
rect 265 92 269 96
rect 271 92 275 96
rect 277 92 281 96
rect 343 92 347 96
rect 349 92 353 96
rect 355 92 359 96
rect 361 92 365 96
rect 367 92 371 96
rect 433 92 437 96
rect 439 92 443 96
rect 445 92 449 96
rect 451 92 455 96
rect 457 92 461 96
rect 523 92 527 96
rect 529 92 533 96
rect 535 92 539 96
rect 541 92 545 96
rect 547 92 551 96
rect 613 92 617 96
rect 619 92 623 96
rect 625 92 629 96
rect 631 92 635 96
rect 637 92 641 96
rect 703 92 707 96
rect 709 92 713 96
rect 715 92 719 96
rect 721 92 725 96
rect 727 92 731 96
rect 793 92 797 96
rect 799 92 803 96
rect 805 92 809 96
rect 811 92 815 96
rect 817 92 821 96
rect 883 92 887 96
rect 889 92 893 96
rect 895 92 899 96
rect 901 92 905 96
rect 907 92 911 96
rect 973 92 977 96
rect 979 92 983 96
rect 985 92 989 96
rect 991 92 995 96
rect 997 92 1001 96
rect 1063 92 1067 96
rect 1069 92 1073 96
rect 1075 92 1079 96
rect 1081 92 1085 96
rect 1087 92 1091 96
rect 1153 92 1157 96
rect 1159 92 1163 96
rect 1165 92 1169 96
rect 1171 92 1175 96
rect 1177 92 1181 96
rect 1243 92 1247 96
rect 1249 92 1253 96
rect 1255 92 1259 96
rect 1261 92 1265 96
rect 1267 92 1271 96
rect 1333 92 1337 96
rect 1339 92 1343 96
rect 1345 92 1349 96
rect 1351 92 1355 96
rect 1357 92 1361 96
<< psubstratepcontact >>
rect 122 1373 126 1377
rect 123 1364 127 1368
rect 131 1364 135 1368
<< nsubstratencontact >>
rect 136 1414 140 1418
rect 153 1415 157 1419
rect 128 1410 132 1414
<< pad >>
rect 142 1454 212 1524
rect 232 1454 302 1524
rect 322 1454 392 1524
rect 412 1454 482 1524
rect 502 1454 572 1524
rect 592 1454 662 1524
rect 682 1454 752 1524
rect 772 1454 842 1524
rect 862 1454 932 1524
rect 952 1454 1022 1524
rect 1042 1454 1112 1524
rect 1132 1454 1202 1524
rect 1222 1454 1292 1524
rect 1312 1454 1382 1524
rect 0 1312 70 1382
rect 1454 1312 1524 1382
rect 0 1222 70 1292
rect 1454 1222 1524 1292
rect 0 1132 70 1202
rect 1454 1132 1524 1202
rect 0 1042 70 1112
rect 1454 1042 1524 1112
rect 0 952 70 1022
rect 1454 952 1524 1022
rect 0 862 70 932
rect 1454 862 1524 932
rect 0 772 70 842
rect 1454 772 1524 842
rect 0 682 70 752
rect 1454 682 1524 752
rect 0 592 70 662
rect 1454 592 1524 662
rect 0 502 70 572
rect 1454 502 1524 572
rect 0 412 70 482
rect 1454 412 1524 482
rect 0 322 70 392
rect 1454 322 1524 392
rect 0 232 70 302
rect 1454 232 1524 302
rect 0 142 70 212
rect 1454 142 1524 212
rect 142 0 212 70
rect 232 0 302 70
rect 322 0 392 70
rect 412 0 482 70
rect 502 0 572 70
rect 592 0 662 70
rect 682 0 752 70
rect 772 0 842 70
rect 862 0 932 70
rect 952 0 1022 70
rect 1042 0 1112 70
rect 1132 0 1202 70
rect 1222 0 1292 70
rect 1312 0 1382 70
<< glass >>
rect 0 1488 1524 1524
rect 0 1485 356 1488
rect 359 1485 1524 1488
rect 0 1454 1524 1485
rect 0 70 70 1454
rect 1454 70 1524 1454
rect 0 0 1524 70
use Porta_CMOS_part1  Porta_CMOS_part1_0
timestamp 1609148708
transform 1 0 126 0 1 1402
box -4 -19 8 6
use Porta_CMOS_part2  Porta_CMOS_part2_0
timestamp 1609157506
transform 1 0 154 0 1 1401
box -12 -35 16 11
<< labels >>
rlabel pad 27 1345 27 1345 1 vA!
rlabel pad 31 1260 31 1260 1 vB!
rlabel pad 33 1163 33 1163 1 vC!
rlabel pad 178 1489 178 1489 1 Vdd!
rlabel pad 1347 34 1347 34 1 GND!
rlabel pad 265 1493 265 1493 1 vF!
<< end >>
