Practica 2 simulació de l'inversor resposta dinamica (Tasca 5)
.include mosfet.model
*.include inversorCMOS.spice

*Capacitat residual dels transistors
*CL 3 0 1p

vi 1 0 0 pulse(0 5V 0s 1fs 1fs 10ns 20ns)
Vdd 2 0 5V
Mn 3 1 0 0 nfet W=3u L=2u
Mp 3 1 2 2 pfet W=3u L=2u


.tran 20p 200ns 0 20p
*.tran printMostresAlTerminal tempsFinal tempsInical SeparacioEntreMostres

*.dc vinput 0 5 0.1 
.control
run
plot v(1) v(3)
plot -i(vdd)
.endc
.end