magic
tech scmos
timestamp 1605178259
<< nwell >>
rect -3 15 11 41
<< polysilicon >>
rect -2 25 2 27
rect 5 25 7 27
rect -2 5 0 25
rect -2 3 2 5
rect 5 3 7 5
<< ndiffusion >>
rect 2 5 5 6
rect 2 2 5 3
<< pdiffusion >>
rect 2 27 5 28
rect 2 24 5 25
<< metal1 >>
rect -8 37 2 41
rect 6 37 20 41
rect -8 32 20 37
rect 2 17 6 20
rect -12 12 -6 16
rect 2 14 15 17
rect 2 10 6 14
rect -9 -2 2 2
rect 6 -2 13 2
rect 17 -2 18 2
rect -9 -7 18 -2
<< ntransistor >>
rect 2 3 5 5
<< ptransistor >>
rect 2 25 5 27
<< polycontact >>
rect -6 12 -2 16
<< ndcontact >>
rect 2 6 6 10
rect 2 -2 6 2
<< pdcontact >>
rect 2 28 6 32
rect 2 20 6 24
<< psubstratepcontact >>
rect 13 -2 17 2
<< nsubstratencontact >>
rect 2 37 6 41
<< labels >>
rlabel metal1 -6 34 -6 34 1 Vdd!
rlabel metal1 14 15 14 15 1 Vo
rlabel metal1 -11 14 -11 14 3 Vi
rlabel metal1 -7 -3 -7 -3 2 Gnd!
<< end >>
