magic
tech scmos
timestamp 1608810559
<< nwell >>
rect -4 -5 9 8
<< polysilicon >>
rect 1 1 4 3
rect 7 1 9 3
rect 1 -8 3 1
rect -4 -10 3 -8
rect 1 -19 3 -10
rect 1 -21 4 -19
rect 7 -21 9 -19
<< ndiffusion >>
rect 4 -19 7 -18
rect 4 -22 7 -21
<< pdiffusion >>
rect 4 3 7 4
rect 4 0 7 1
<< metal1 >>
rect 0 5 4 8
rect 8 5 9 8
rect 4 -7 8 -4
rect 4 -11 9 -7
rect 4 -14 8 -11
rect 0 -26 4 -23
rect 8 -26 9 -23
<< ntransistor >>
rect 4 -21 7 -19
<< ptransistor >>
rect 4 1 7 3
<< ndcontact >>
rect 4 -18 8 -14
rect 4 -26 8 -22
<< pdcontact >>
rect 4 4 8 8
rect 4 -4 8 0
<< psubstratepcontact >>
rect -4 -26 0 -22
<< nsubstratencontact >>
rect -4 4 0 8
<< labels >>
rlabel metal1 1 6 1 6 5 Vdd!
rlabel metal1 1 -25 1 -25 1 GND!
rlabel polysilicon -3 -9 -3 -9 3 vA!
rlabel metal1 7 -9 7 -9 7 vnA!
<< end >>
