Practica 2 simulació de l'inversor (Tasca 4)
.include mosfet.model
.include inversorCMOS.spice

*Extracció
vinput Vi Gnd dc 0

*Font d'alimentacio
Vddfont Vdd Gnd dc 5

.dc vinput 0 5 0.1
.control
run
plot v(vo)
plot -i(vddfont)
.endc
.end