magic
tech scmos
timestamp 1609157506
<< nwell >>
rect -12 -15 16 11
<< polysilicon >>
rect -5 9 -3 11
rect 1 9 3 11
rect 6 9 8 11
rect -5 -5 -3 -4
rect -8 -6 -3 -5
rect -10 -7 -3 -6
rect -12 -8 -6 -7
rect -12 -9 -8 -8
rect -12 -19 -10 -9
rect -12 -21 -6 -19
rect -8 -23 -5 -21
rect -7 -25 -5 -23
rect 1 -25 3 -15
rect 6 -17 8 -15
rect 6 -19 11 -17
rect 9 -25 11 -19
rect -7 -35 -5 -33
rect 1 -35 3 -33
rect 9 -35 11 -33
<< ndiffusion >>
rect -8 -33 -7 -25
rect -5 -33 -4 -25
rect 0 -33 1 -25
rect 3 -29 4 -25
rect 8 -29 9 -25
rect 3 -33 9 -29
rect 11 -33 12 -25
<< pdiffusion >>
rect -6 -4 -5 9
rect -3 -4 1 9
rect -2 -8 1 -4
rect 0 -15 1 -8
rect 3 -15 6 9
rect 8 -12 9 9
rect 8 -15 12 -12
<< metal1 >>
rect -12 9 16 11
rect -12 -4 -10 9
rect -6 7 9 9
rect 13 -12 16 9
rect -4 -19 0 -15
rect -3 -22 16 -19
rect 4 -25 8 -22
rect -12 -35 -8 -33
rect 0 -33 12 -32
rect -4 -35 16 -33
<< ntransistor >>
rect -7 -33 -5 -25
rect 1 -33 3 -25
rect 9 -33 11 -25
<< ptransistor >>
rect -5 -4 -3 9
rect 1 -15 3 9
rect 6 -15 8 9
<< ndcontact >>
rect -12 -33 -8 -25
rect -4 -33 0 -25
rect 4 -29 8 -25
rect 12 -33 16 -25
<< pdcontact >>
rect -10 -4 -6 9
rect -4 -15 0 -8
rect 9 -12 13 9
<< labels >>
rlabel metal1 -10 7 -10 7 4 Vdd!
rlabel polysilicon 2 -19 2 -19 1 vB!
rlabel polysilicon 7 -19 7 -19 1 vC!
rlabel polysilicon -10 -20 -10 -20 3 vnA!
rlabel metal1 13 -20 13 -20 7 vF!
rlabel metal1 -10 -34 -10 -34 2 GND!
<< end >>
